module fpu_mul( clk, rst, enable, opa, opb, sign, product_7, exponent_5);
input		clk;
input		rst;
input		enable;
input	[63:0]	opa, opb;
output		sign;
output  [55:0] product_7;
output  [11:0] exponent_5;

reg [5:0] 	product_shift;
reg [5:0] 	product_shift_2;


reg   sign;
reg   [51:0] mantissa_a;
reg   [51:0] mantissa_b;
reg   [10:0] exponent_a;
reg   [10:0] exponent_b;
reg		a_is_norm;
reg		b_is_norm;
reg		a_is_zero; 
reg		b_is_zero; 
reg		in_zero;
reg   [11:0] exponent_terms;
reg    exponent_gt_expoffset;
reg   [11:0] exponent_under;
reg   [11:0] exponent_1;
wire   [11:0] exponent = 0;
reg   [11:0] exponent_2;
reg   exponent_gt_prodshift;
reg   [11:0] exponent_3;
reg   [11:0] exponent_4;
reg  exponent_et_zero;
reg   [52:0] mul_a;
reg   [52:0] mul_b;
reg   [105:0] product;
reg   [105:0] product_1;
reg   [105:0] product_2;
reg   [105:0] product_3;
reg   [105:0] product_4; 
reg   [105:0] product_5;
reg   [105:0] product_6;
reg		product_lsb; // if there are any 1's in the remainder
wire  [55:0] product_7 =  { 1'b0, product_6[105:52], product_lsb }; 
reg  [11:0] exponent_5;		
task booth_final;
    input [52:0] in1, in2;
    output [105:0] out;
    begin
      q = in1;
      m = in2;
      q1 = 1'b0;
      acc = 52'b0;
      count = 53;

      if (count > 0) begin
        for (count = 53; count > 0; count = count - 1) begin
          check = {q[0], q1};
          if (check == 2'b00 || check == 2'b11) begin
            y = q[0];
            {acc[52:0], q[52:0], q1} = {acc[52:0], q[52:0], q1} >> 1;
            acc[52:0] = {y, acc[51:0]};
          end
          else if (check == 2'b10) begin
            y = q[0];
            y1 = ~m + 1'b1;
            acc = acc + y1;
            {acc[52:0], q[52:0], q1} = {acc[52:0], q[52:0], q1} >> 1;
            acc[52:0] = {y, acc[51:0]};
          end
          else begin
            y = q[0];
            acc = acc + m;
            {acc[52:0], q[52:0], q1} = {acc[52:0], q[52:0], q1} >> 1;
            acc[52:0] = {y, acc[51:0]};
          end
        end
        out = {acc, q};
      end
      else
        out = {acc, q};
    end
 endtask
always @(posedge clk) 
begin
	if (rst) begin
		sign <= 0;
		mantissa_a <= 0;
		mantissa_b <= 0;
		exponent_a <= 0;
		exponent_b <= 0;
		a_is_norm <= 0;
		b_is_norm <= 0;
		a_is_zero <= 0; 
		b_is_zero <= 0; 
		in_zero <= 0;
		exponent_terms <= 0;
		exponent_gt_expoffset <= 0;
		exponent_under <= 0;
		exponent_1 <= 0; 
		exponent_2 <= 0;
		exponent_gt_prodshift <= 0;
		exponent_3 <= 0;
		exponent_4 <= 0;
		exponent_et_zero <= 0;
		mul_a <= 0; 
		mul_b <= 0;
		product <= 0;
		product_1 <= 0;
		product_2 <= 0; 
		product_3 <= 0;
		product_4 <= 0;
		product_5 <= 0; 
		product_6 <= 0;
		product_lsb <= 0;
		exponent_5 <= 0;
		product_shift_2 <= 0;
	end
	else if (enable) begin
		sign <= opa[63] ^ opb[63];
		mantissa_a <= opa[51:0];
		mantissa_b <= opb[51:0];
		exponent_a <= opa[62:52];
		exponent_b <= opb[62:52];
		a_is_norm <= |exponent_a;
		b_is_norm <= |exponent_b;
		a_is_zero <= !(|opa[62:0]); 
		b_is_zero <= !(|opb[62:0]); 
		in_zero <= a_is_zero | b_is_zero;
		exponent_terms <= exponent_a + exponent_b + !a_is_norm + !b_is_norm;
		exponent_gt_expoffset <= exponent_terms > 1021;
		exponent_under <= 1022 - exponent_terms;
		exponent_1 <= exponent_terms - 1022; 
		exponent_2 <= exponent_gt_expoffset ? exponent_1 : exponent;
		exponent_gt_prodshift <= exponent_2 > product_shift_2;
		exponent_3 <= exponent_2 - product_shift;
		exponent_4 <= exponent_gt_prodshift ? exponent_3 : exponent;
		exponent_et_zero <= exponent_4 == 0;
		mul_a <= { a_is_norm, mantissa_a };
		mul_b <= { b_is_norm, mantissa_b };
		booth_final(mul_a,mul_b,product) //calling and using task
		product_1 <= product >> exponent_under;
		product_2 <= exponent_gt_expoffset ? product : product_1; 
		product_3 <= product_2 << product_shift_2;
		product_4 <= product_2 << exponent_2;
		product_5 <= exponent_gt_prodshift ? product_3  : product_4;
		product_6 <= exponent_et_zero ? product_5 >> 1 : product_5;
		product_lsb <= |product_6[51:0];
		exponent_5 <= in_zero ? 12'b0 : exponent_4;
		product_shift_2 <= product_shift; // redundant register
			// reduces fanout on product_shift
	end
end

always @(product)
   casex(product)	
    106'b1?????????????????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  0;
	106'b01????????????????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  1;
	106'b001???????????????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  2;
	106'b0001??????????????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  3;
	106'b00001?????????????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  4;
	106'b000001????????????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  5;
	106'b0000001???????????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  6;
	106'b00000001??????????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  7;
	106'b000000001?????????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  8;
	106'b0000000001????????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  9;
	106'b00000000001???????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  10;
	106'b000000000001??????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  11;
	106'b0000000000001?????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  12;
	106'b00000000000001????????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  13;
	106'b000000000000001???????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  14;
	106'b0000000000000001??????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  15;
	106'b00000000000000001?????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  16;
	106'b000000000000000001????????????????????????????????????????????????????????????????????????????????????????: product_shift <=  17;
	106'b0000000000000000001???????????????????????????????????????????????????????????????????????????????????????: product_shift <=  18;
	106'b00000000000000000001??????????????????????????????????????????????????????????????????????????????????????: product_shift <=  19;
	106'b000000000000000000001?????????????????????????????????????????????????????????????????????????????????????: product_shift <=  20;
	106'b0000000000000000000001????????????????????????????????????????????????????????????????????????????????????: product_shift <=  21;
	106'b00000000000000000000001???????????????????????????????????????????????????????????????????????????????????: product_shift <=  22;
	106'b000000000000000000000001??????????????????????????????????????????????????????????????????????????????????: product_shift <=  23;
	106'b0000000000000000000000001?????????????????????????????????????????????????????????????????????????????????: product_shift <=  24;
	106'b00000000000000000000000001????????????????????????????????????????????????????????????????????????????????: product_shift <=  25;
	106'b000000000000000000000000001???????????????????????????????????????????????????????????????????????????????: product_shift <=  26;
	106'b0000000000000000000000000001??????????????????????????????????????????????????????????????????????????????: product_shift <=  27;
	106'b00000000000000000000000000001?????????????????????????????????????????????????????????????????????????????: product_shift <=  28;
	106'b000000000000000000000000000001????????????????????????????????????????????????????????????????????????????: product_shift <=  29;
	106'b0000000000000000000000000000001???????????????????????????????????????????????????????????????????????????: product_shift <=  30;
	106'b00000000000000000000000000000001??????????????????????????????????????????????????????????????????????????: product_shift <=  31;
	106'b000000000000000000000000000000001?????????????????????????????????????????????????????????????????????????: product_shift <=  32;
	106'b0000000000000000000000000000000001????????????????????????????????????????????????????????????????????????: product_shift <=  33;
	106'b00000000000000000000000000000000001???????????????????????????????????????????????????????????????????????: product_shift <=  34;
	106'b000000000000000000000000000000000001??????????????????????????????????????????????????????????????????????: product_shift <=  35;
	106'b0000000000000000000000000000000000001?????????????????????????????????????????????????????????????????????: product_shift <=  36;
	106'b00000000000000000000000000000000000001????????????????????????????????????????????????????????????????????: product_shift <=  37;
	106'b000000000000000000000000000000000000001???????????????????????????????????????????????????????????????????: product_shift <=  38;
	106'b0000000000000000000000000000000000000001??????????????????????????????????????????????????????????????????: product_shift <=  39;
	106'b00000000000000000000000000000000000000001?????????????????????????????????????????????????????????????????: product_shift <=  40;
	106'b000000000000000000000000000000000000000001????????????????????????????????????????????????????????????????: product_shift <=  41;
	106'b0000000000000000000000000000000000000000001???????????????????????????????????????????????????????????????: product_shift <=  42;
	106'b00000000000000000000000000000000000000000001??????????????????????????????????????????????????????????????: product_shift <=  43;
	106'b000000000000000000000000000000000000000000001?????????????????????????????????????????????????????????????: product_shift <=  44;
	106'b0000000000000000000000000000000000000000000001????????????????????????????????????????????????????????????: product_shift <=  45;
	106'b00000000000000000000000000000000000000000000001???????????????????????????????????????????????????????????: product_shift <=  46;
	106'b000000000000000000000000000000000000000000000001??????????????????????????????????????????????????????????: product_shift <=  47;
	106'b0000000000000000000000000000000000000000000000001?????????????????????????????????????????????????????????: product_shift <=  48;
    106'b00000000000000000000000000000000000000000000000001????????????????????????????????????????????????????????: product_shift <=  49;
	106'b000000000000000000000000000000000000000000000000001???????????????????????????????????????????????????????: product_shift <=  50;
	106'b0000000000000000000000000000000000000000000000000001??????????????????????????????????????????????????????: product_shift <=  51;
	106'b00000000000000000000000000000000000000000000000000001?????????????????????????????????????????????????????: product_shift <=  52;
	106'b000000000000000000000000000000000000000000000000000000????????????????????????????????????????????????????: product_shift <=  53;
	  // It's not necessary to go past 53, because you will only get more than 53 zeros
	  // when multiplying 2 denormalized numbers together, in which case you will underflow
	endcase	

endmodule
